class Transaction;

// stimulus 
rand 